`timescale 1ns/1ns
//Part 1:
module MUX_4x1(input a,b,c,d, input [1:0] S, output f);
 assign #(36,38) f = S[1] ? (S[0] ? d : c) : (S[0] ? b : a);
endmodule

//Part 2:
module Barrel_shifter_4bit(input [1:0] N, input [3:0] A, output [3:0] SHO);
 MUX_4x1 MUX1(A[0],A[1],A[2],A[3], N, SHO[0]), MUX2(A[1],A[2],A[3],A[0], N, SHO[1]),
         MUX3(A[2],A[3],A[0],A[1], N, SHO[2]), MUX4(A[3],A[0],A[1],A[2], N, SHO[3]);
endmodule

//Part 3:
module MUX_16x1(input [15:0] I, input [3:0] S, output f);
reg [3:0] w;
 MUX_4x1 MUX1(I[0],I[1],I[2],I[3], {S[1],S[0]}, w[0]),
         MUX2(I[4],I[5],I[6],I[7], {S[1],S[0]}, w[1]),
         MUX3(I[8],I[9],I[10],I[11], {S[1],S[0]}, w[2]),
         MUX4(I[12],I[13],I[14],I[15], {S[1],S[0]}, w[3]),
         MUX5(w[0],w[1],w[2],w[3], {S[3],S[2]}, f);
endmodule

//Part 4:
module Barrel_shifter_16x1(input [15:0] I, input [3:0] S, output [15:0] SHO);
MUX_16x1 MUX1({I[15],I[14],I[13],I[12],I[11],I[10],I[9],I[8],I[7],I[6],I[5],I[4],I[3],I[2],I[1],I[0]},S,SHO[0]),
         MUX2({I[0],I[15],I[14],I[13],I[12],I[11],I[10],I[9],I[8],I[7],I[6],I[5],I[4],I[3],I[2],I[1]},S,SHO[1]),
         MUX3({I[1],I[0],I[15],I[14],I[13],I[12],I[11],I[10],I[9],I[8],I[7],I[6],I[5],I[4],I[3],I[2]},S,SHO[2]),
         MUX4({I[2],I[1],I[0],I[15],I[14],I[13],I[12],I[11],I[10],I[9],I[8],I[7],I[6],I[5],I[4],I[3]},S,SHO[3]),
         MUX5({I[3],I[2],I[1],I[0],I[15],I[14],I[13],I[12],I[11],I[10],I[9],I[8],I[7],I[6],I[5],I[4]},S,SHO[4]),
         MUX6({I[4],I[3],I[2],I[1],I[0],I[15],I[14],I[13],I[12],I[11],I[10],I[9],I[8],I[7],I[6],I[5]},S,SHO[5]),
         MUX7({I[5],I[4],I[3],I[2],I[1],I[0],I[15],I[14],I[13],I[12],I[11],I[10],I[9],I[8],I[7],I[6]},S,SHO[6]),
         MUX8({I[6],I[5],I[4],I[3],I[2],I[1],I[0],I[15],I[14],I[13],I[12],I[11],I[10],I[9],I[8],I[7]},S,SHO[7]),
         MUX9({I[7],I[6],I[5],I[4],I[3],I[2],I[1],I[0],I[15],I[14],I[13],I[12],I[11],I[10],I[9],I[8]},S,SHO[8]),
         MUX10({I[8],I[7],I[6],I[5],I[4],I[3],I[2],I[1],I[0],I[15],I[14],I[13],I[12],I[11],I[10],I[9]},S,SHO[9]),
         MUX11({I[9],I[8],I[7],I[6],I[5],I[4],I[3],I[2],I[1],I[0],I[15],I[14],I[13],I[12],I[11],I[10]},S,SHO[10]),
         MUX12({I[10],I[9],I[8],I[7],I[6],I[5],I[4],I[3],I[2],I[1],I[0],I[15],I[14],I[13],I[12],I[11]},S,SHO[11]),
         MUX13({I[11],I[10],I[9],I[8],I[7],I[6],I[5],I[4],I[3],I[2],I[1],I[0],I[15],I[14],I[13],I[12]},S,SHO[12]),
         MUX14({I[12],I[11],I[10],I[9],I[8],I[7],I[6],I[5],I[4],I[3],I[2],I[1],I[0],I[15],I[14],I[13]},S,SHO[13]),
         MUX15({I[13],I[12],I[11],I[10],I[9],I[8],I[7],I[6],I[5],I[4],I[3],I[2],I[1],I[0],I[15],I[14]},S,SHO[14]),
         MUX16({I[14],I[13],I[12],I[11],I[10],I[9],I[8],I[7],I[6],I[5],I[4],I[3],I[2],I[1],I[0],I[15]},S,SHO[15]);
endmodule